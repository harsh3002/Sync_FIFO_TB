`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"